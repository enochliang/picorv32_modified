module fi_wrapper;
//=============================
// Tasks
//=============================

task setmask;
  input [31:0] num;
  output [63:0] o_mask;
  begin
    o_mask = 1 << num;
  end
endtask

task cycle2num;
  input [31:0] cyc;
  output [55:0] num;
  begin
    num2char(cyc/1000000,num[55:48]);
    cyc = cyc % 1000000;
    num2char(cyc/100000,num[47:40]);
    cyc = cyc % 100000;
    num2char(cyc/10000,num[39:32]);
    cyc = cyc % 10000;
    num2char(cyc/1000,num[31:24]);
    cyc = cyc % 1000;
    num2char(cyc/100,num[23:16]);
    cyc = cyc % 100;
    num2char(cyc/10,num[15:8]);
    cyc = cyc % 10;

    num2char(cyc,num[7:0]);
  end
endtask

task num2char;
  input [31:0] num;
  output [7:0] ch;
  begin
    case(num)
      'd0:ch=8'd48;
      'd1:ch=8'd49;
      'd2:ch=8'd50;
      'd3:ch=8'd51;
      'd4:ch=8'd52;
      'd5:ch=8'd53;
      'd6:ch=8'd54;
      'd7:ch=8'd55;
      'd8:ch=8'd56;
      'd9:ch=8'd57;
    endcase
  end
endtask

task num2str;
  input [31:0] num;
  output [31:0] str;
  begin
    num2char(num/1000,str[31:24]);
    num = num % 1000;
    num2char(num/100,str[23:16]);
    num = num % 100;
    num2char(num/10,str[15:8]);
    num = num % 10;

    num2char(num,str[7:0]);
  end
endtask
//----------------------------------------------------------------
//  FI_Wrapper Control Signals Declaration
//----------------------------------------------------------------
reg tb_clk;
reg [31:0] cycle;
reg [55:0] cycle_str;
reg [55:0] cycle_str2;
reg [31:0] inj_id;
reg [31:0] inj_id_str;
reg [31:0] bit_pos;
reg [31:0] bit_pos_str;
reg [63:0] mask;
reg inj_flag;
reg input_flag;
//=====================
// input port buffers
//=====================
reg [0:0] tb_in__resetn;
reg [0:0] tb_in2__resetn;
reg [0:0] tb_in__mem_axi_awready;
reg [0:0] tb_in2__mem_axi_awready;
reg [0:0] tb_in__mem_axi_wready;
reg [0:0] tb_in2__mem_axi_wready;
reg [0:0] tb_in__mem_axi_bvalid;
reg [0:0] tb_in2__mem_axi_bvalid;
reg [0:0] tb_in__mem_axi_arready;
reg [0:0] tb_in2__mem_axi_arready;
reg [0:0] tb_in__mem_axi_rvalid;
reg [0:0] tb_in2__mem_axi_rvalid;
reg [31:0] tb_in__mem_axi_rdata;
reg [31:0] tb_in2__mem_axi_rdata;
reg [0:0] tb_in__pcpi_wr;
reg [0:0] tb_in2__pcpi_wr;
reg [31:0] tb_in__pcpi_rd;
reg [31:0] tb_in2__pcpi_rd;
reg [0:0] tb_in__pcpi_wait;
reg [0:0] tb_in2__pcpi_wait;
reg [0:0] tb_in__pcpi_ready;
reg [0:0] tb_in2__pcpi_ready;
reg [31:0] tb_in__irq;
reg [31:0] tb_in2__irq;
//=====================
// output port buffers
//=====================
reg [0:0] tb_out__trap;
reg [0:0] tb_out__mem_axi_awvalid;
reg [31:0] tb_out__mem_axi_awaddr;
reg [0:0] tb_out__mem_axi_wvalid;
reg [31:0] tb_out__mem_axi_wdata;
reg [3:0] tb_out__mem_axi_wstrb;
reg [0:0] tb_out__mem_axi_bready;
reg [0:0] tb_out__mem_axi_arvalid;
reg [31:0] tb_out__mem_axi_araddr;
reg [2:0] tb_out__mem_axi_arprot;
reg [0:0] tb_out__mem_axi_rready;
reg [0:0] tb_out__pcpi_valid;
reg [31:0] tb_out__pcpi_insn;
reg [31:0] tb_out__pcpi_rs1;
reg [31:0] tb_out__pcpi_rs2;
reg [31:0] tb_out__eoi;
reg [0:0] tb_out__trace_valid;
reg [35:0] tb_out__trace_data;
//=====================
// output port wire
//=====================
wire [0:0] trap;
wire [0:0] mem_axi_awvalid;
wire [31:0] mem_axi_awaddr;
wire [0:0] mem_axi_wvalid;
wire [31:0] mem_axi_wdata;
wire [3:0] mem_axi_wstrb;
wire [0:0] mem_axi_bready;
wire [0:0] mem_axi_arvalid;
wire [31:0] mem_axi_araddr;
wire [2:0] mem_axi_arprot;
wire [0:0] mem_axi_rready;
wire [0:0] pcpi_valid;
wire [31:0] pcpi_insn;
wire [31:0] pcpi_rs1;
wire [31:0] pcpi_rs2;
wire [31:0] eoi;
wire [0:0] trace_valid;
wire [35:0] trace_data;
//=============================
// fault free register buffers
//=============================
reg [0:0] ff_buf__picorv32_axi__axi_adapter__ack_awvalid;
reg [0:0] ff_buf__picorv32_axi__axi_adapter__ack_arvalid;
reg [0:0] ff_buf__picorv32_axi__axi_adapter__ack_wvalid;
reg [0:0] ff_buf__picorv32_axi__axi_adapter__xfer_done;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__trap_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_valid_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_instr_reg;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__mem_addr_reg;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__mem_wdata_reg;
reg [3:0] ff_buf__picorv32_axi__picorv32_core__mem_wstrb_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__pcpi_valid_reg;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__pcpi_insn_reg;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__eoi_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__trace_valid_reg;
reg [35:0] ff_buf__picorv32_axi__picorv32_core__trace_data_reg;
reg [63:0] ff_buf__picorv32_axi__picorv32_core__count_cycle;
reg [63:0] ff_buf__picorv32_axi__picorv32_core__count_instr;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__reg_pc;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__reg_next_pc;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__reg_op1;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__reg_op2;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__reg_out;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__reg_sh;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__next_insn_opcode;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__dbg_insn_addr;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__irq_delay;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__irq_active;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__irq_mask;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__irq_pending;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__timer;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__0;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__1;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__2;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__3;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__4;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__5;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__6;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__7;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__8;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__9;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__10;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__11;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__12;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__13;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__14;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__15;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__16;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__17;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__18;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__19;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__20;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__21;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__22;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__23;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__24;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__25;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__26;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__27;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__28;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__29;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__30;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__31;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__32;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__33;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__34;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cpuregs__35;
reg [1:0] ff_buf__picorv32_axi__picorv32_core__mem_state;
reg [1:0] ff_buf__picorv32_axi__picorv32_core__mem_wordsize;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__mem_rdata_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_do_prefetch;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_do_rinst;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_do_rdata;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_do_wdata;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_la_secondword;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__mem_la_firstword_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__last_mem_valid;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__prefetched_high_word;
reg [15:0] ff_buf__picorv32_axi__picorv32_core__mem_16bit_buffer;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_lui;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_auipc;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_jal;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_jalr;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_beq;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_bne;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_blt;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_bge;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_bltu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_bgeu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_lb;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_lh;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_lw;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_lbu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_lhu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sb;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sh;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sw;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_addi;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_slti;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sltiu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_xori;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_ori;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_andi;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_slli;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_srli;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_srai;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_add;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sub;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sll;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_slt;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sltu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_xor;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_srl;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_sra;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_or;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_and;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_rdcycle;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_rdcycleh;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_rdinstr;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_rdinstrh;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_ecall_ebreak;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_fence;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_getq;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_setq;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_retirq;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_maskirq;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_waitirq;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__instr_timer;
reg [5:0] ff_buf__picorv32_axi__picorv32_core__decoded_rd;
reg [5:0] ff_buf__picorv32_axi__picorv32_core__decoded_rs1;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__decoded_rs2;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__decoded_imm;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__decoded_imm_j;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__decoder_trigger;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__decoder_trigger_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__compressed_instr;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_lb_lh_lw_lbu_lhu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_slli_srli_srai;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_jalr_addi_slti_sltiu_xori_ori_andi;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_sb_sh_sw;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_sll_srl_sra;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal_jalr_addi_add_sub;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_slti_blt_slt;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_sltiu_bltu_sltu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_beq_bne_blt_bge_bltu_bgeu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_lbu_lhu_lw;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_alu_reg_imm;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_alu_reg_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__is_compare;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__dbg_rs1val;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__dbg_rs2val;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__dbg_rs1val_valid;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__dbg_rs2val_valid;
reg [63:0] ff_buf__picorv32_axi__picorv32_core__q_ascii_instr;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__q_insn_imm;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__q_insn_opcode;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__q_insn_rs1;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__q_insn_rs2;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__q_insn_rd;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__dbg_next;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__dbg_valid_insn;
reg [63:0] ff_buf__picorv32_axi__picorv32_core__cached_ascii_instr;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cached_insn_imm;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__cached_insn_opcode;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__cached_insn_rs1;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__cached_insn_rs2;
reg [4:0] ff_buf__picorv32_axi__picorv32_core__cached_insn_rd;
reg [7:0] ff_buf__picorv32_axi__picorv32_core__cpu_state;
reg [1:0] ff_buf__picorv32_axi__picorv32_core__irq_state;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_store;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_stalu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_branch;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_compr;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_trace;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_is_lu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_is_lh;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__latched_is_lb;
reg [5:0] ff_buf__picorv32_axi__picorv32_core__latched_rd;
reg [3:0] ff_buf__picorv32_axi__picorv32_core__pcpi_timeout_counter;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__pcpi_timeout;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__do_waitirq;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__alu_out_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__alu_out_0_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__alu_wait;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__alu_wait_2;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__clear_prefetched_high_word_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__shift_out;
reg [3:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__active;
reg [32:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1;
reg [32:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2;
reg [32:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1_q;
reg [32:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2_q;
reg [63:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd;
reg [63:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__pcpi_insn_valid_q;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wr_reg;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_rd_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_ready_reg;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_div;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_divu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_rem;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_remu;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_q;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__dividend;
reg [62:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__divisor;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient;
reg [31:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient_msk;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__running;
reg [0:0] ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__outsign;
//=============================
// golden register buffers
//=============================
reg [0:0] golden_buf__picorv32_axi__axi_adapter__ack_awvalid;
reg [0:0] golden_buf__picorv32_axi__axi_adapter__ack_arvalid;
reg [0:0] golden_buf__picorv32_axi__axi_adapter__ack_wvalid;
reg [0:0] golden_buf__picorv32_axi__axi_adapter__xfer_done;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__trap_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_valid_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_instr_reg;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__mem_addr_reg;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__mem_wdata_reg;
reg [3:0] golden_buf__picorv32_axi__picorv32_core__mem_wstrb_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__pcpi_valid_reg;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__pcpi_insn_reg;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__eoi_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__trace_valid_reg;
reg [35:0] golden_buf__picorv32_axi__picorv32_core__trace_data_reg;
reg [63:0] golden_buf__picorv32_axi__picorv32_core__count_cycle;
reg [63:0] golden_buf__picorv32_axi__picorv32_core__count_instr;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__reg_pc;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__reg_next_pc;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__reg_op1;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__reg_op2;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__reg_out;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__reg_sh;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__next_insn_opcode;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__dbg_insn_addr;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__irq_delay;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__irq_active;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__irq_mask;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__irq_pending;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__timer;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__0;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__1;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__2;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__3;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__4;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__5;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__6;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__7;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__8;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__9;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__10;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__11;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__12;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__13;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__14;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__15;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__16;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__17;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__18;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__19;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__20;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__21;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__22;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__23;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__24;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__25;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__26;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__27;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__28;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__29;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__30;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__31;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__32;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__33;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__34;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cpuregs__35;
reg [1:0] golden_buf__picorv32_axi__picorv32_core__mem_state;
reg [1:0] golden_buf__picorv32_axi__picorv32_core__mem_wordsize;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__mem_rdata_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_do_prefetch;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_do_rinst;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_do_rdata;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_do_wdata;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_la_secondword;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__mem_la_firstword_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__last_mem_valid;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__prefetched_high_word;
reg [15:0] golden_buf__picorv32_axi__picorv32_core__mem_16bit_buffer;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_lui;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_auipc;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_jal;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_jalr;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_beq;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_bne;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_blt;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_bge;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_bltu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_bgeu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_lb;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_lh;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_lw;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_lbu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_lhu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sb;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sh;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sw;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_addi;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_slti;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sltiu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_xori;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_ori;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_andi;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_slli;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_srli;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_srai;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_add;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sub;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sll;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_slt;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sltu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_xor;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_srl;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_sra;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_or;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_and;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_rdcycle;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_rdcycleh;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_rdinstr;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_rdinstrh;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_ecall_ebreak;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_fence;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_getq;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_setq;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_retirq;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_maskirq;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_waitirq;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__instr_timer;
reg [5:0] golden_buf__picorv32_axi__picorv32_core__decoded_rd;
reg [5:0] golden_buf__picorv32_axi__picorv32_core__decoded_rs1;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__decoded_rs2;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__decoded_imm;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__decoded_imm_j;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__decoder_trigger;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__decoder_trigger_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__compressed_instr;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_lb_lh_lw_lbu_lhu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_slli_srli_srai;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_jalr_addi_slti_sltiu_xori_ori_andi;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_sb_sh_sw;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_sll_srl_sra;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal_jalr_addi_add_sub;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_slti_blt_slt;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_sltiu_bltu_sltu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_beq_bne_blt_bge_bltu_bgeu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_lbu_lhu_lw;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_alu_reg_imm;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_alu_reg_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__is_compare;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__dbg_rs1val;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__dbg_rs2val;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__dbg_rs1val_valid;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__dbg_rs2val_valid;
reg [63:0] golden_buf__picorv32_axi__picorv32_core__q_ascii_instr;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__q_insn_imm;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__q_insn_opcode;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__q_insn_rs1;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__q_insn_rs2;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__q_insn_rd;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__dbg_next;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__dbg_valid_insn;
reg [63:0] golden_buf__picorv32_axi__picorv32_core__cached_ascii_instr;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cached_insn_imm;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__cached_insn_opcode;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__cached_insn_rs1;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__cached_insn_rs2;
reg [4:0] golden_buf__picorv32_axi__picorv32_core__cached_insn_rd;
reg [7:0] golden_buf__picorv32_axi__picorv32_core__cpu_state;
reg [1:0] golden_buf__picorv32_axi__picorv32_core__irq_state;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_store;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_stalu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_branch;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_compr;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_trace;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_is_lu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_is_lh;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__latched_is_lb;
reg [5:0] golden_buf__picorv32_axi__picorv32_core__latched_rd;
reg [3:0] golden_buf__picorv32_axi__picorv32_core__pcpi_timeout_counter;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__pcpi_timeout;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__do_waitirq;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__alu_out_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__alu_out_0_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__alu_wait;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__alu_wait_2;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__clear_prefetched_high_word_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__shift_out;
reg [3:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__active;
reg [32:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1;
reg [32:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2;
reg [32:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1_q;
reg [32:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2_q;
reg [63:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd;
reg [63:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__pcpi_insn_valid_q;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wr_reg;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_rd_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_ready_reg;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_div;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_divu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_rem;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_remu;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_q;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__dividend;
reg [62:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__divisor;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient;
reg [31:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient_msk;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__running;
reg [0:0] golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__outsign;


	picorv32_axi #(
		.COMPRESSED_ISA(1),
		.ENABLE_FAST_MUL(1),
		.ENABLE_DIV(1),
		.ENABLE_IRQ(1),
		.ENABLE_TRACE(1)
	) picorv32_axi (
	    .clk(tb_clk),
            .resetn(tb_in__resetn),
            .mem_axi_awready(tb_in__mem_axi_awready),
            .mem_axi_wready(tb_in__mem_axi_wready),
            .mem_axi_bvalid(tb_in__mem_axi_bvalid),
            .mem_axi_arready(tb_in__mem_axi_arready),
            .mem_axi_rvalid(tb_in__mem_axi_rvalid),
            .mem_axi_rdata(tb_in__mem_axi_rdata),
            .pcpi_wr(tb_in__pcpi_wr),
            .pcpi_rd(tb_in__pcpi_rd),
            .pcpi_wait(tb_in__pcpi_wait),
            .pcpi_ready(tb_in__pcpi_ready),
            .irq(tb_in__irq),
            .trap(trap),
            .mem_axi_awvalid(mem_axi_awvalid),
            .mem_axi_awaddr(mem_axi_awaddr),
            .mem_axi_wvalid(mem_axi_wvalid),
            .mem_axi_wdata(mem_axi_wdata),
            .mem_axi_wstrb(mem_axi_wstrb),
            .mem_axi_bready(mem_axi_bready),
            .mem_axi_arvalid(mem_axi_arvalid),
            .mem_axi_araddr(mem_axi_araddr),
            .mem_axi_arprot(mem_axi_arprot),
            .mem_axi_rready(mem_axi_rready),
            .pcpi_valid(pcpi_valid),
            .pcpi_insn(pcpi_insn),
            .pcpi_rs1(pcpi_rs1),
            .pcpi_rs2(pcpi_rs2),
            .eoi(eoi),
            .trace_valid(trace_valid),
            .trace_data(trace_data),
          );

// File IO
integer f_control,f_input,f_golden,f_observe;
initial begin
  tb_clk = 0;
  inj_flag = 0;
  input_flag = 0;

  f_control = $fopen("control.txt","r");
  $fscanf(f_control, "%d", cycle);
  $fscanf(f_control, "%d", inj_id);
  $fscanf(f_control, "%d", bit_pos);
  $fclose(f_control);

  num2str(inj_id, inj_id_str);
  num2str(bit_pos, bit_pos_str);
  cycle2num(cycle,cycle_str);
  cycle2num(cycle+1,cycle_str2);
  setmask(bit_pos, mask);

  //==============================
  // load fault free input buffer
  //==============================
  f_input = $fopen({"ff_value/ff_value_C",cycle_str,".txt"},"r");
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__axi_adapter__ack_awvalid);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__axi_adapter__ack_arvalid);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__axi_adapter__ack_wvalid);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__axi_adapter__xfer_done);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__trap_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_valid_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_instr_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_addr_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_wdata_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_wstrb_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__pcpi_valid_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__pcpi_insn_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__eoi_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__trace_valid_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__trace_data_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__count_cycle);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__count_instr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__reg_pc);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__reg_next_pc);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__reg_op1);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__reg_op2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__reg_out);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__reg_sh);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__next_insn_opcode);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_insn_addr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__irq_delay);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__irq_active);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__irq_mask);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__irq_pending);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__timer);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__0);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__1);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__3);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__4);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__5);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__6);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__7);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__8);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__9);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__10);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__11);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__12);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__13);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__14);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__15);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__16);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__17);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__18);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__19);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__20);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__21);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__22);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__23);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__24);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__25);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__26);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__27);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__28);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__29);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__30);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__31);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__32);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__33);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__34);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpuregs__35);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_state);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_wordsize);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_rdata_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_do_prefetch);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_do_rinst);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_do_rdata);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_do_wdata);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_la_secondword);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_la_firstword_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__last_mem_valid);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__prefetched_high_word);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__mem_16bit_buffer);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_lui);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_auipc);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_jal);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_jalr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_beq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_bne);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_blt);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_bge);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_bltu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_bgeu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_lb);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_lh);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_lw);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_lbu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_lhu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sb);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sh);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sw);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_addi);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_slti);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sltiu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_xori);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_ori);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_andi);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_slli);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_srli);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_srai);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_add);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sub);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sll);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_slt);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sltu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_xor);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_srl);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_sra);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_or);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_and);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_rdcycle);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_rdcycleh);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_rdinstr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_rdinstrh);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_ecall_ebreak);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_fence);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_getq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_setq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_retirq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_maskirq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_waitirq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__instr_timer);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoded_rd);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoded_rs1);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoded_rs2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoded_imm);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoded_imm_j);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoder_trigger);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoder_trigger_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__compressed_instr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_lb_lh_lw_lbu_lhu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_slli_srli_srai);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_jalr_addi_slti_sltiu_xori_ori_andi);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_sb_sh_sw);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_sll_srl_sra);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal_jalr_addi_add_sub);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_slti_blt_slt);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_sltiu_bltu_sltu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_beq_bne_blt_bge_bltu_bgeu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_lbu_lhu_lw);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_alu_reg_imm);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_alu_reg_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__is_compare);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_rs1val);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_rs2val);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_rs1val_valid);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_rs2val_valid);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__q_ascii_instr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__q_insn_imm);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__q_insn_opcode);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__q_insn_rs1);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__q_insn_rs2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__q_insn_rd);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_next);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__dbg_valid_insn);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cached_ascii_instr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cached_insn_imm);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cached_insn_opcode);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cached_insn_rs1);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cached_insn_rs2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cached_insn_rd);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__cpu_state);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__irq_state);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_store);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_stalu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_branch);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_compr);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_trace);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_is_lu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_is_lh);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_is_lb);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__latched_rd);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__pcpi_timeout_counter);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__pcpi_timeout);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__do_waitirq);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__alu_out_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__alu_out_0_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__alu_wait);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__alu_wait_2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__clear_prefetched_high_word_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__shift_out);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__active);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__pcpi_insn_valid_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wr_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_rd_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_ready_reg);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_div);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_divu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_rem);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_remu);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_q);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__dividend);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__divisor);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient_msk);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__running);
  $fscanf(f_input,"%b",ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__outsign);
  $fscanf(f_input,"%b",tb_in__resetn);
  $fscanf(f_input,"%b",tb_in__mem_axi_awready);
  $fscanf(f_input,"%b",tb_in__mem_axi_wready);
  $fscanf(f_input,"%b",tb_in__mem_axi_bvalid);
  $fscanf(f_input,"%b",tb_in__mem_axi_arready);
  $fscanf(f_input,"%b",tb_in__mem_axi_rvalid);
  $fscanf(f_input,"%b",tb_in__mem_axi_rdata);
  $fscanf(f_input,"%b",tb_in__pcpi_wr);
  $fscanf(f_input,"%b",tb_in__pcpi_rd);
  $fscanf(f_input,"%b",tb_in__pcpi_wait);
  $fscanf(f_input,"%b",tb_in__pcpi_ready);
  $fscanf(f_input,"%b",tb_in__irq);
  $fscanf(f_input,"%b",tb_in2__resetn);
  $fscanf(f_input,"%b",tb_in2__mem_axi_awready);
  $fscanf(f_input,"%b",tb_in2__mem_axi_wready);
  $fscanf(f_input,"%b",tb_in2__mem_axi_bvalid);
  $fscanf(f_input,"%b",tb_in2__mem_axi_arready);
  $fscanf(f_input,"%b",tb_in2__mem_axi_rvalid);
  $fscanf(f_input,"%b",tb_in2__mem_axi_rdata);
  $fscanf(f_input,"%b",tb_in2__pcpi_wr);
  $fscanf(f_input,"%b",tb_in2__pcpi_rd);
  $fscanf(f_input,"%b",tb_in2__pcpi_wait);
  $fscanf(f_input,"%b",tb_in2__pcpi_ready);
  $fscanf(f_input,"%b",tb_in2__irq);
  //==============================
  // load golden output buffer
  //==============================
  f_golden = $fopen({"golden_value/golden_value_C",cycle_str2,".txt"},"r");
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__axi_adapter__ack_awvalid);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__axi_adapter__ack_arvalid);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__axi_adapter__ack_wvalid);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__axi_adapter__xfer_done);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__trap_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_valid_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_instr_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_addr_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_wdata_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_wstrb_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__pcpi_valid_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__pcpi_insn_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__eoi_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__trace_valid_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__trace_data_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__count_cycle);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__count_instr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__reg_pc);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__reg_next_pc);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__reg_op1);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__reg_op2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__reg_out);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__reg_sh);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__next_insn_opcode);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_insn_addr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__irq_delay);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__irq_active);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__irq_mask);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__irq_pending);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__timer);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__0);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__1);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__3);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__4);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__5);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__6);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__7);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__8);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__9);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__10);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__11);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__12);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__13);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__14);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__15);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__16);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__17);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__18);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__19);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__20);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__21);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__22);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__23);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__24);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__25);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__26);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__27);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__28);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__29);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__30);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__31);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__32);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__33);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__34);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpuregs__35);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_state);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_wordsize);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_rdata_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_do_prefetch);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_do_rinst);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_do_rdata);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_do_wdata);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_la_secondword);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_la_firstword_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__last_mem_valid);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__prefetched_high_word);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__mem_16bit_buffer);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_lui);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_auipc);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_jal);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_jalr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_beq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_bne);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_blt);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_bge);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_bltu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_bgeu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_lb);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_lh);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_lw);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_lbu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_lhu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sb);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sh);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sw);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_addi);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_slti);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sltiu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_xori);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_ori);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_andi);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_slli);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_srli);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_srai);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_add);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sub);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sll);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_slt);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sltu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_xor);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_srl);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_sra);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_or);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_and);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_rdcycle);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_rdcycleh);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_rdinstr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_rdinstrh);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_ecall_ebreak);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_fence);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_getq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_setq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_retirq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_maskirq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_waitirq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__instr_timer);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoded_rd);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoded_rs1);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoded_rs2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoded_imm);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoded_imm_j);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoder_trigger);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoder_trigger_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__compressed_instr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_lb_lh_lw_lbu_lhu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_slli_srli_srai);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_jalr_addi_slti_sltiu_xori_ori_andi);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_sb_sh_sw);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_sll_srl_sra);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal_jalr_addi_add_sub);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_slti_blt_slt);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_sltiu_bltu_sltu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_beq_bne_blt_bge_bltu_bgeu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_lbu_lhu_lw);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_alu_reg_imm);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_alu_reg_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__is_compare);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_rs1val);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_rs2val);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_rs1val_valid);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_rs2val_valid);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__q_ascii_instr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__q_insn_imm);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__q_insn_opcode);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__q_insn_rs1);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__q_insn_rs2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__q_insn_rd);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_next);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__dbg_valid_insn);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cached_ascii_instr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cached_insn_imm);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cached_insn_opcode);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cached_insn_rs1);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cached_insn_rs2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cached_insn_rd);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__cpu_state);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__irq_state);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_store);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_stalu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_branch);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_compr);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_trace);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_is_lu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_is_lh);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_is_lb);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__latched_rd);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__pcpi_timeout_counter);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__pcpi_timeout);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__do_waitirq);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__alu_out_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__alu_out_0_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__alu_wait);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__alu_wait_2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__clear_prefetched_high_word_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__shift_out);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__active);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__pcpi_insn_valid_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wr_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_rd_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_ready_reg);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_div);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_divu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_rem);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_remu);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_q);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__dividend);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__divisor);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient_msk);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__running);
  $fscanf(f_golden,"%b",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__outsign);
  //================
  // timing control
  //================
  #CLK_HALF_PERIOD input_flag = !input_flag;
  #CLK_HALF_PERIOD inj_flag = !inj_flag;
  #CLK_HALF_PERIOD tb_clk = !tb_clk;
  #CLK_HALF_PERIOD input_flag = !input_flag;
  #CLK_HALF_PERIOD tb_clk = !tb_clk;
  #CLK_HALF_PERIOD;
  //===============================
  // dump fault effect observation
  //===============================
  f_observe = $fopen({"result/result_C", cycle_str, "_R", inj_id_str, "_B", pos_bit_str , ".txt"},"r");
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__axi_adapter__ack_awvalid^picorv32_axi.axi_adapter.ack_awvalid);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__axi_adapter__ack_arvalid^picorv32_axi.axi_adapter.ack_arvalid);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__axi_adapter__ack_wvalid^picorv32_axi.axi_adapter.ack_wvalid);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__axi_adapter__xfer_done^picorv32_axi.axi_adapter.xfer_done);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__trap_reg^picorv32_axi.picorv32_core.trap_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_valid_reg^picorv32_axi.picorv32_core.mem_valid_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_instr_reg^picorv32_axi.picorv32_core.mem_instr_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_addr_reg^picorv32_axi.picorv32_core.mem_addr_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_wdata_reg^picorv32_axi.picorv32_core.mem_wdata_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_wstrb_reg^picorv32_axi.picorv32_core.mem_wstrb_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__pcpi_valid_reg^picorv32_axi.picorv32_core.pcpi_valid_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__pcpi_insn_reg^picorv32_axi.picorv32_core.pcpi_insn_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__eoi_reg^picorv32_axi.picorv32_core.eoi_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__trace_valid_reg^picorv32_axi.picorv32_core.trace_valid_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__trace_data_reg^picorv32_axi.picorv32_core.trace_data_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__count_cycle^picorv32_axi.picorv32_core.count_cycle);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__count_instr^picorv32_axi.picorv32_core.count_instr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__reg_pc^picorv32_axi.picorv32_core.reg_pc);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__reg_next_pc^picorv32_axi.picorv32_core.reg_next_pc);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__reg_op1^picorv32_axi.picorv32_core.reg_op1);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__reg_op2^picorv32_axi.picorv32_core.reg_op2);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__reg_out^picorv32_axi.picorv32_core.reg_out);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__reg_sh^picorv32_axi.picorv32_core.reg_sh);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__next_insn_opcode^picorv32_axi.picorv32_core.next_insn_opcode);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_insn_addr^picorv32_axi.picorv32_core.dbg_insn_addr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__irq_delay^picorv32_axi.picorv32_core.irq_delay);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__irq_active^picorv32_axi.picorv32_core.irq_active);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__irq_mask^picorv32_axi.picorv32_core.irq_mask);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__irq_pending^picorv32_axi.picorv32_core.irq_pending);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__timer^picorv32_axi.picorv32_core.timer);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__0^picorv32_axi.picorv32_core.cpuregs[0]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__1^picorv32_axi.picorv32_core.cpuregs[1]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__2^picorv32_axi.picorv32_core.cpuregs[2]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__3^picorv32_axi.picorv32_core.cpuregs[3]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__4^picorv32_axi.picorv32_core.cpuregs[4]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__5^picorv32_axi.picorv32_core.cpuregs[5]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__6^picorv32_axi.picorv32_core.cpuregs[6]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__7^picorv32_axi.picorv32_core.cpuregs[7]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__8^picorv32_axi.picorv32_core.cpuregs[8]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__9^picorv32_axi.picorv32_core.cpuregs[9]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__10^picorv32_axi.picorv32_core.cpuregs[10]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__11^picorv32_axi.picorv32_core.cpuregs[11]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__12^picorv32_axi.picorv32_core.cpuregs[12]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__13^picorv32_axi.picorv32_core.cpuregs[13]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__14^picorv32_axi.picorv32_core.cpuregs[14]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__15^picorv32_axi.picorv32_core.cpuregs[15]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__16^picorv32_axi.picorv32_core.cpuregs[16]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__17^picorv32_axi.picorv32_core.cpuregs[17]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__18^picorv32_axi.picorv32_core.cpuregs[18]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__19^picorv32_axi.picorv32_core.cpuregs[19]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__20^picorv32_axi.picorv32_core.cpuregs[20]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__21^picorv32_axi.picorv32_core.cpuregs[21]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__22^picorv32_axi.picorv32_core.cpuregs[22]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__23^picorv32_axi.picorv32_core.cpuregs[23]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__24^picorv32_axi.picorv32_core.cpuregs[24]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__25^picorv32_axi.picorv32_core.cpuregs[25]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__26^picorv32_axi.picorv32_core.cpuregs[26]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__27^picorv32_axi.picorv32_core.cpuregs[27]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__28^picorv32_axi.picorv32_core.cpuregs[28]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__29^picorv32_axi.picorv32_core.cpuregs[29]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__30^picorv32_axi.picorv32_core.cpuregs[30]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__31^picorv32_axi.picorv32_core.cpuregs[31]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__32^picorv32_axi.picorv32_core.cpuregs[32]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__33^picorv32_axi.picorv32_core.cpuregs[33]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__34^picorv32_axi.picorv32_core.cpuregs[34]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpuregs__35^picorv32_axi.picorv32_core.cpuregs[35]);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_state^picorv32_axi.picorv32_core.mem_state);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_wordsize^picorv32_axi.picorv32_core.mem_wordsize);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_rdata_q^picorv32_axi.picorv32_core.mem_rdata_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_do_prefetch^picorv32_axi.picorv32_core.mem_do_prefetch);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_do_rinst^picorv32_axi.picorv32_core.mem_do_rinst);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_do_rdata^picorv32_axi.picorv32_core.mem_do_rdata);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_do_wdata^picorv32_axi.picorv32_core.mem_do_wdata);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_la_secondword^picorv32_axi.picorv32_core.mem_la_secondword);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_la_firstword_reg^picorv32_axi.picorv32_core.mem_la_firstword_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__last_mem_valid^picorv32_axi.picorv32_core.last_mem_valid);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__prefetched_high_word^picorv32_axi.picorv32_core.prefetched_high_word);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__mem_16bit_buffer^picorv32_axi.picorv32_core.mem_16bit_buffer);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_lui^picorv32_axi.picorv32_core.instr_lui);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_auipc^picorv32_axi.picorv32_core.instr_auipc);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_jal^picorv32_axi.picorv32_core.instr_jal);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_jalr^picorv32_axi.picorv32_core.instr_jalr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_beq^picorv32_axi.picorv32_core.instr_beq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_bne^picorv32_axi.picorv32_core.instr_bne);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_blt^picorv32_axi.picorv32_core.instr_blt);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_bge^picorv32_axi.picorv32_core.instr_bge);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_bltu^picorv32_axi.picorv32_core.instr_bltu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_bgeu^picorv32_axi.picorv32_core.instr_bgeu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_lb^picorv32_axi.picorv32_core.instr_lb);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_lh^picorv32_axi.picorv32_core.instr_lh);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_lw^picorv32_axi.picorv32_core.instr_lw);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_lbu^picorv32_axi.picorv32_core.instr_lbu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_lhu^picorv32_axi.picorv32_core.instr_lhu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sb^picorv32_axi.picorv32_core.instr_sb);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sh^picorv32_axi.picorv32_core.instr_sh);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sw^picorv32_axi.picorv32_core.instr_sw);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_addi^picorv32_axi.picorv32_core.instr_addi);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_slti^picorv32_axi.picorv32_core.instr_slti);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sltiu^picorv32_axi.picorv32_core.instr_sltiu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_xori^picorv32_axi.picorv32_core.instr_xori);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_ori^picorv32_axi.picorv32_core.instr_ori);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_andi^picorv32_axi.picorv32_core.instr_andi);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_slli^picorv32_axi.picorv32_core.instr_slli);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_srli^picorv32_axi.picorv32_core.instr_srli);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_srai^picorv32_axi.picorv32_core.instr_srai);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_add^picorv32_axi.picorv32_core.instr_add);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sub^picorv32_axi.picorv32_core.instr_sub);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sll^picorv32_axi.picorv32_core.instr_sll);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_slt^picorv32_axi.picorv32_core.instr_slt);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sltu^picorv32_axi.picorv32_core.instr_sltu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_xor^picorv32_axi.picorv32_core.instr_xor);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_srl^picorv32_axi.picorv32_core.instr_srl);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_sra^picorv32_axi.picorv32_core.instr_sra);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_or^picorv32_axi.picorv32_core.instr_or);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_and^picorv32_axi.picorv32_core.instr_and);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_rdcycle^picorv32_axi.picorv32_core.instr_rdcycle);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_rdcycleh^picorv32_axi.picorv32_core.instr_rdcycleh);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_rdinstr^picorv32_axi.picorv32_core.instr_rdinstr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_rdinstrh^picorv32_axi.picorv32_core.instr_rdinstrh);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_ecall_ebreak^picorv32_axi.picorv32_core.instr_ecall_ebreak);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_fence^picorv32_axi.picorv32_core.instr_fence);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_getq^picorv32_axi.picorv32_core.instr_getq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_setq^picorv32_axi.picorv32_core.instr_setq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_retirq^picorv32_axi.picorv32_core.instr_retirq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_maskirq^picorv32_axi.picorv32_core.instr_maskirq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_waitirq^picorv32_axi.picorv32_core.instr_waitirq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__instr_timer^picorv32_axi.picorv32_core.instr_timer);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoded_rd^picorv32_axi.picorv32_core.decoded_rd);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoded_rs1^picorv32_axi.picorv32_core.decoded_rs1);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoded_rs2^picorv32_axi.picorv32_core.decoded_rs2);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoded_imm^picorv32_axi.picorv32_core.decoded_imm);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoded_imm_j^picorv32_axi.picorv32_core.decoded_imm_j);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoder_trigger^picorv32_axi.picorv32_core.decoder_trigger);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoder_trigger_q^picorv32_axi.picorv32_core.decoder_trigger_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger^picorv32_axi.picorv32_core.decoder_pseudo_trigger);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger_q^picorv32_axi.picorv32_core.decoder_pseudo_trigger_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__compressed_instr^picorv32_axi.picorv32_core.compressed_instr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal^picorv32_axi.picorv32_core.is_lui_auipc_jal);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_lb_lh_lw_lbu_lhu^picorv32_axi.picorv32_core.is_lb_lh_lw_lbu_lhu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_slli_srli_srai^picorv32_axi.picorv32_core.is_slli_srli_srai);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_jalr_addi_slti_sltiu_xori_ori_andi^picorv32_axi.picorv32_core.is_jalr_addi_slti_sltiu_xori_ori_andi);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_sb_sh_sw^picorv32_axi.picorv32_core.is_sb_sh_sw);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_sll_srl_sra^picorv32_axi.picorv32_core.is_sll_srl_sra);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal_jalr_addi_add_sub^picorv32_axi.picorv32_core.is_lui_auipc_jal_jalr_addi_add_sub);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_slti_blt_slt^picorv32_axi.picorv32_core.is_slti_blt_slt);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_sltiu_bltu_sltu^picorv32_axi.picorv32_core.is_sltiu_bltu_sltu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_beq_bne_blt_bge_bltu_bgeu^picorv32_axi.picorv32_core.is_beq_bne_blt_bge_bltu_bgeu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_lbu_lhu_lw^picorv32_axi.picorv32_core.is_lbu_lhu_lw);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_alu_reg_imm^picorv32_axi.picorv32_core.is_alu_reg_imm);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_alu_reg_reg^picorv32_axi.picorv32_core.is_alu_reg_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__is_compare^picorv32_axi.picorv32_core.is_compare);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_rs1val^picorv32_axi.picorv32_core.dbg_rs1val);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_rs2val^picorv32_axi.picorv32_core.dbg_rs2val);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_rs1val_valid^picorv32_axi.picorv32_core.dbg_rs1val_valid);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_rs2val_valid^picorv32_axi.picorv32_core.dbg_rs2val_valid);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__q_ascii_instr^picorv32_axi.picorv32_core.q_ascii_instr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__q_insn_imm^picorv32_axi.picorv32_core.q_insn_imm);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__q_insn_opcode^picorv32_axi.picorv32_core.q_insn_opcode);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__q_insn_rs1^picorv32_axi.picorv32_core.q_insn_rs1);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__q_insn_rs2^picorv32_axi.picorv32_core.q_insn_rs2);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__q_insn_rd^picorv32_axi.picorv32_core.q_insn_rd);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_next^picorv32_axi.picorv32_core.dbg_next);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__dbg_valid_insn^picorv32_axi.picorv32_core.dbg_valid_insn);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cached_ascii_instr^picorv32_axi.picorv32_core.cached_ascii_instr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cached_insn_imm^picorv32_axi.picorv32_core.cached_insn_imm);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cached_insn_opcode^picorv32_axi.picorv32_core.cached_insn_opcode);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cached_insn_rs1^picorv32_axi.picorv32_core.cached_insn_rs1);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cached_insn_rs2^picorv32_axi.picorv32_core.cached_insn_rs2);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cached_insn_rd^picorv32_axi.picorv32_core.cached_insn_rd);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__cpu_state^picorv32_axi.picorv32_core.cpu_state);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__irq_state^picorv32_axi.picorv32_core.irq_state);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_store^picorv32_axi.picorv32_core.latched_store);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_stalu^picorv32_axi.picorv32_core.latched_stalu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_branch^picorv32_axi.picorv32_core.latched_branch);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_compr^picorv32_axi.picorv32_core.latched_compr);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_trace^picorv32_axi.picorv32_core.latched_trace);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_is_lu^picorv32_axi.picorv32_core.latched_is_lu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_is_lh^picorv32_axi.picorv32_core.latched_is_lh);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_is_lb^picorv32_axi.picorv32_core.latched_is_lb);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__latched_rd^picorv32_axi.picorv32_core.latched_rd);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__pcpi_timeout_counter^picorv32_axi.picorv32_core.pcpi_timeout_counter);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__pcpi_timeout^picorv32_axi.picorv32_core.pcpi_timeout);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__do_waitirq^picorv32_axi.picorv32_core.do_waitirq);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__alu_out_q^picorv32_axi.picorv32_core.alu_out_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__alu_out_0_q^picorv32_axi.picorv32_core.alu_out_0_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__alu_wait^picorv32_axi.picorv32_core.alu_wait);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__alu_wait_2^picorv32_axi.picorv32_core.alu_wait_2);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__clear_prefetched_high_word_q^picorv32_axi.picorv32_core.clear_prefetched_high_word_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__shift_out^picorv32_axi.picorv32_core.genblk1.pcpi_mul.shift_out);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__active^picorv32_axi.picorv32_core.genblk1.pcpi_mul.active);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1^picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2^picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1_q^picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2_q^picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd^picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd_q^picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__pcpi_insn_valid_q^picorv32_axi.picorv32_core.genblk1.pcpi_mul.pcpi_insn_valid_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wr_reg^picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wr_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_rd_reg^picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_rd_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_reg^picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_ready_reg^picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_ready_reg);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_div^picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_div);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_divu^picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_divu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_rem^picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_rem);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_remu^picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_remu);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_q^picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_q);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__dividend^picorv32_axi.picorv32_core.genblk2.pcpi_div.dividend);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__divisor^picorv32_axi.picorv32_core.genblk2.pcpi_div.divisor);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient^picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient_msk^picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient_msk);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__running^picorv32_axi.picorv32_core.genblk2.pcpi_div.running);
  $fwrite(f_observe,"%b\n",golden_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__outsign^picorv32_axi.picorv32_core.genblk2.pcpi_div.outsign);
end
//===============================
// always blocks
//===============================
// fault free pattern filling (to registers)
always@(posedge input_flag)begin
  picorv32_axi.axi_adapter.ack_awvalid <= ff_buf__picorv32_axi__axi_adapter__ack_awvalid;
  picorv32_axi.axi_adapter.ack_arvalid <= ff_buf__picorv32_axi__axi_adapter__ack_arvalid;
  picorv32_axi.axi_adapter.ack_wvalid <= ff_buf__picorv32_axi__axi_adapter__ack_wvalid;
  picorv32_axi.axi_adapter.xfer_done <= ff_buf__picorv32_axi__axi_adapter__xfer_done;
  picorv32_axi.picorv32_core.trap_reg <= ff_buf__picorv32_axi__picorv32_core__trap_reg;
  picorv32_axi.picorv32_core.mem_valid_reg <= ff_buf__picorv32_axi__picorv32_core__mem_valid_reg;
  picorv32_axi.picorv32_core.mem_instr_reg <= ff_buf__picorv32_axi__picorv32_core__mem_instr_reg;
  picorv32_axi.picorv32_core.mem_addr_reg <= ff_buf__picorv32_axi__picorv32_core__mem_addr_reg;
  picorv32_axi.picorv32_core.mem_wdata_reg <= ff_buf__picorv32_axi__picorv32_core__mem_wdata_reg;
  picorv32_axi.picorv32_core.mem_wstrb_reg <= ff_buf__picorv32_axi__picorv32_core__mem_wstrb_reg;
  picorv32_axi.picorv32_core.pcpi_valid_reg <= ff_buf__picorv32_axi__picorv32_core__pcpi_valid_reg;
  picorv32_axi.picorv32_core.pcpi_insn_reg <= ff_buf__picorv32_axi__picorv32_core__pcpi_insn_reg;
  picorv32_axi.picorv32_core.eoi_reg <= ff_buf__picorv32_axi__picorv32_core__eoi_reg;
  picorv32_axi.picorv32_core.trace_valid_reg <= ff_buf__picorv32_axi__picorv32_core__trace_valid_reg;
  picorv32_axi.picorv32_core.trace_data_reg <= ff_buf__picorv32_axi__picorv32_core__trace_data_reg;
  picorv32_axi.picorv32_core.count_cycle <= ff_buf__picorv32_axi__picorv32_core__count_cycle;
  picorv32_axi.picorv32_core.count_instr <= ff_buf__picorv32_axi__picorv32_core__count_instr;
  picorv32_axi.picorv32_core.reg_pc <= ff_buf__picorv32_axi__picorv32_core__reg_pc;
  picorv32_axi.picorv32_core.reg_next_pc <= ff_buf__picorv32_axi__picorv32_core__reg_next_pc;
  picorv32_axi.picorv32_core.reg_op1 <= ff_buf__picorv32_axi__picorv32_core__reg_op1;
  picorv32_axi.picorv32_core.reg_op2 <= ff_buf__picorv32_axi__picorv32_core__reg_op2;
  picorv32_axi.picorv32_core.reg_out <= ff_buf__picorv32_axi__picorv32_core__reg_out;
  picorv32_axi.picorv32_core.reg_sh <= ff_buf__picorv32_axi__picorv32_core__reg_sh;
  picorv32_axi.picorv32_core.next_insn_opcode <= ff_buf__picorv32_axi__picorv32_core__next_insn_opcode;
  picorv32_axi.picorv32_core.dbg_insn_addr <= ff_buf__picorv32_axi__picorv32_core__dbg_insn_addr;
  picorv32_axi.picorv32_core.irq_delay <= ff_buf__picorv32_axi__picorv32_core__irq_delay;
  picorv32_axi.picorv32_core.irq_active <= ff_buf__picorv32_axi__picorv32_core__irq_active;
  picorv32_axi.picorv32_core.irq_mask <= ff_buf__picorv32_axi__picorv32_core__irq_mask;
  picorv32_axi.picorv32_core.irq_pending <= ff_buf__picorv32_axi__picorv32_core__irq_pending;
  picorv32_axi.picorv32_core.timer <= ff_buf__picorv32_axi__picorv32_core__timer;
  picorv32_axi.picorv32_core.cpuregs[0] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__0;
  picorv32_axi.picorv32_core.cpuregs[1] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__1;
  picorv32_axi.picorv32_core.cpuregs[2] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__2;
  picorv32_axi.picorv32_core.cpuregs[3] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__3;
  picorv32_axi.picorv32_core.cpuregs[4] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__4;
  picorv32_axi.picorv32_core.cpuregs[5] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__5;
  picorv32_axi.picorv32_core.cpuregs[6] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__6;
  picorv32_axi.picorv32_core.cpuregs[7] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__7;
  picorv32_axi.picorv32_core.cpuregs[8] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__8;
  picorv32_axi.picorv32_core.cpuregs[9] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__9;
  picorv32_axi.picorv32_core.cpuregs[10] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__10;
  picorv32_axi.picorv32_core.cpuregs[11] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__11;
  picorv32_axi.picorv32_core.cpuregs[12] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__12;
  picorv32_axi.picorv32_core.cpuregs[13] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__13;
  picorv32_axi.picorv32_core.cpuregs[14] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__14;
  picorv32_axi.picorv32_core.cpuregs[15] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__15;
  picorv32_axi.picorv32_core.cpuregs[16] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__16;
  picorv32_axi.picorv32_core.cpuregs[17] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__17;
  picorv32_axi.picorv32_core.cpuregs[18] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__18;
  picorv32_axi.picorv32_core.cpuregs[19] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__19;
  picorv32_axi.picorv32_core.cpuregs[20] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__20;
  picorv32_axi.picorv32_core.cpuregs[21] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__21;
  picorv32_axi.picorv32_core.cpuregs[22] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__22;
  picorv32_axi.picorv32_core.cpuregs[23] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__23;
  picorv32_axi.picorv32_core.cpuregs[24] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__24;
  picorv32_axi.picorv32_core.cpuregs[25] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__25;
  picorv32_axi.picorv32_core.cpuregs[26] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__26;
  picorv32_axi.picorv32_core.cpuregs[27] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__27;
  picorv32_axi.picorv32_core.cpuregs[28] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__28;
  picorv32_axi.picorv32_core.cpuregs[29] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__29;
  picorv32_axi.picorv32_core.cpuregs[30] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__30;
  picorv32_axi.picorv32_core.cpuregs[31] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__31;
  picorv32_axi.picorv32_core.cpuregs[32] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__32;
  picorv32_axi.picorv32_core.cpuregs[33] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__33;
  picorv32_axi.picorv32_core.cpuregs[34] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__34;
  picorv32_axi.picorv32_core.cpuregs[35] <= ff_buf__picorv32_axi__picorv32_core__cpuregs__35;
  picorv32_axi.picorv32_core.mem_state <= ff_buf__picorv32_axi__picorv32_core__mem_state;
  picorv32_axi.picorv32_core.mem_wordsize <= ff_buf__picorv32_axi__picorv32_core__mem_wordsize;
  picorv32_axi.picorv32_core.mem_rdata_q <= ff_buf__picorv32_axi__picorv32_core__mem_rdata_q;
  picorv32_axi.picorv32_core.mem_do_prefetch <= ff_buf__picorv32_axi__picorv32_core__mem_do_prefetch;
  picorv32_axi.picorv32_core.mem_do_rinst <= ff_buf__picorv32_axi__picorv32_core__mem_do_rinst;
  picorv32_axi.picorv32_core.mem_do_rdata <= ff_buf__picorv32_axi__picorv32_core__mem_do_rdata;
  picorv32_axi.picorv32_core.mem_do_wdata <= ff_buf__picorv32_axi__picorv32_core__mem_do_wdata;
  picorv32_axi.picorv32_core.mem_la_secondword <= ff_buf__picorv32_axi__picorv32_core__mem_la_secondword;
  picorv32_axi.picorv32_core.mem_la_firstword_reg <= ff_buf__picorv32_axi__picorv32_core__mem_la_firstword_reg;
  picorv32_axi.picorv32_core.last_mem_valid <= ff_buf__picorv32_axi__picorv32_core__last_mem_valid;
  picorv32_axi.picorv32_core.prefetched_high_word <= ff_buf__picorv32_axi__picorv32_core__prefetched_high_word;
  picorv32_axi.picorv32_core.mem_16bit_buffer <= ff_buf__picorv32_axi__picorv32_core__mem_16bit_buffer;
  picorv32_axi.picorv32_core.instr_lui <= ff_buf__picorv32_axi__picorv32_core__instr_lui;
  picorv32_axi.picorv32_core.instr_auipc <= ff_buf__picorv32_axi__picorv32_core__instr_auipc;
  picorv32_axi.picorv32_core.instr_jal <= ff_buf__picorv32_axi__picorv32_core__instr_jal;
  picorv32_axi.picorv32_core.instr_jalr <= ff_buf__picorv32_axi__picorv32_core__instr_jalr;
  picorv32_axi.picorv32_core.instr_beq <= ff_buf__picorv32_axi__picorv32_core__instr_beq;
  picorv32_axi.picorv32_core.instr_bne <= ff_buf__picorv32_axi__picorv32_core__instr_bne;
  picorv32_axi.picorv32_core.instr_blt <= ff_buf__picorv32_axi__picorv32_core__instr_blt;
  picorv32_axi.picorv32_core.instr_bge <= ff_buf__picorv32_axi__picorv32_core__instr_bge;
  picorv32_axi.picorv32_core.instr_bltu <= ff_buf__picorv32_axi__picorv32_core__instr_bltu;
  picorv32_axi.picorv32_core.instr_bgeu <= ff_buf__picorv32_axi__picorv32_core__instr_bgeu;
  picorv32_axi.picorv32_core.instr_lb <= ff_buf__picorv32_axi__picorv32_core__instr_lb;
  picorv32_axi.picorv32_core.instr_lh <= ff_buf__picorv32_axi__picorv32_core__instr_lh;
  picorv32_axi.picorv32_core.instr_lw <= ff_buf__picorv32_axi__picorv32_core__instr_lw;
  picorv32_axi.picorv32_core.instr_lbu <= ff_buf__picorv32_axi__picorv32_core__instr_lbu;
  picorv32_axi.picorv32_core.instr_lhu <= ff_buf__picorv32_axi__picorv32_core__instr_lhu;
  picorv32_axi.picorv32_core.instr_sb <= ff_buf__picorv32_axi__picorv32_core__instr_sb;
  picorv32_axi.picorv32_core.instr_sh <= ff_buf__picorv32_axi__picorv32_core__instr_sh;
  picorv32_axi.picorv32_core.instr_sw <= ff_buf__picorv32_axi__picorv32_core__instr_sw;
  picorv32_axi.picorv32_core.instr_addi <= ff_buf__picorv32_axi__picorv32_core__instr_addi;
  picorv32_axi.picorv32_core.instr_slti <= ff_buf__picorv32_axi__picorv32_core__instr_slti;
  picorv32_axi.picorv32_core.instr_sltiu <= ff_buf__picorv32_axi__picorv32_core__instr_sltiu;
  picorv32_axi.picorv32_core.instr_xori <= ff_buf__picorv32_axi__picorv32_core__instr_xori;
  picorv32_axi.picorv32_core.instr_ori <= ff_buf__picorv32_axi__picorv32_core__instr_ori;
  picorv32_axi.picorv32_core.instr_andi <= ff_buf__picorv32_axi__picorv32_core__instr_andi;
  picorv32_axi.picorv32_core.instr_slli <= ff_buf__picorv32_axi__picorv32_core__instr_slli;
  picorv32_axi.picorv32_core.instr_srli <= ff_buf__picorv32_axi__picorv32_core__instr_srli;
  picorv32_axi.picorv32_core.instr_srai <= ff_buf__picorv32_axi__picorv32_core__instr_srai;
  picorv32_axi.picorv32_core.instr_add <= ff_buf__picorv32_axi__picorv32_core__instr_add;
  picorv32_axi.picorv32_core.instr_sub <= ff_buf__picorv32_axi__picorv32_core__instr_sub;
  picorv32_axi.picorv32_core.instr_sll <= ff_buf__picorv32_axi__picorv32_core__instr_sll;
  picorv32_axi.picorv32_core.instr_slt <= ff_buf__picorv32_axi__picorv32_core__instr_slt;
  picorv32_axi.picorv32_core.instr_sltu <= ff_buf__picorv32_axi__picorv32_core__instr_sltu;
  picorv32_axi.picorv32_core.instr_xor <= ff_buf__picorv32_axi__picorv32_core__instr_xor;
  picorv32_axi.picorv32_core.instr_srl <= ff_buf__picorv32_axi__picorv32_core__instr_srl;
  picorv32_axi.picorv32_core.instr_sra <= ff_buf__picorv32_axi__picorv32_core__instr_sra;
  picorv32_axi.picorv32_core.instr_or <= ff_buf__picorv32_axi__picorv32_core__instr_or;
  picorv32_axi.picorv32_core.instr_and <= ff_buf__picorv32_axi__picorv32_core__instr_and;
  picorv32_axi.picorv32_core.instr_rdcycle <= ff_buf__picorv32_axi__picorv32_core__instr_rdcycle;
  picorv32_axi.picorv32_core.instr_rdcycleh <= ff_buf__picorv32_axi__picorv32_core__instr_rdcycleh;
  picorv32_axi.picorv32_core.instr_rdinstr <= ff_buf__picorv32_axi__picorv32_core__instr_rdinstr;
  picorv32_axi.picorv32_core.instr_rdinstrh <= ff_buf__picorv32_axi__picorv32_core__instr_rdinstrh;
  picorv32_axi.picorv32_core.instr_ecall_ebreak <= ff_buf__picorv32_axi__picorv32_core__instr_ecall_ebreak;
  picorv32_axi.picorv32_core.instr_fence <= ff_buf__picorv32_axi__picorv32_core__instr_fence;
  picorv32_axi.picorv32_core.instr_getq <= ff_buf__picorv32_axi__picorv32_core__instr_getq;
  picorv32_axi.picorv32_core.instr_setq <= ff_buf__picorv32_axi__picorv32_core__instr_setq;
  picorv32_axi.picorv32_core.instr_retirq <= ff_buf__picorv32_axi__picorv32_core__instr_retirq;
  picorv32_axi.picorv32_core.instr_maskirq <= ff_buf__picorv32_axi__picorv32_core__instr_maskirq;
  picorv32_axi.picorv32_core.instr_waitirq <= ff_buf__picorv32_axi__picorv32_core__instr_waitirq;
  picorv32_axi.picorv32_core.instr_timer <= ff_buf__picorv32_axi__picorv32_core__instr_timer;
  picorv32_axi.picorv32_core.decoded_rd <= ff_buf__picorv32_axi__picorv32_core__decoded_rd;
  picorv32_axi.picorv32_core.decoded_rs1 <= ff_buf__picorv32_axi__picorv32_core__decoded_rs1;
  picorv32_axi.picorv32_core.decoded_rs2 <= ff_buf__picorv32_axi__picorv32_core__decoded_rs2;
  picorv32_axi.picorv32_core.decoded_imm <= ff_buf__picorv32_axi__picorv32_core__decoded_imm;
  picorv32_axi.picorv32_core.decoded_imm_j <= ff_buf__picorv32_axi__picorv32_core__decoded_imm_j;
  picorv32_axi.picorv32_core.decoder_trigger <= ff_buf__picorv32_axi__picorv32_core__decoder_trigger;
  picorv32_axi.picorv32_core.decoder_trigger_q <= ff_buf__picorv32_axi__picorv32_core__decoder_trigger_q;
  picorv32_axi.picorv32_core.decoder_pseudo_trigger <= ff_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger;
  picorv32_axi.picorv32_core.decoder_pseudo_trigger_q <= ff_buf__picorv32_axi__picorv32_core__decoder_pseudo_trigger_q;
  picorv32_axi.picorv32_core.compressed_instr <= ff_buf__picorv32_axi__picorv32_core__compressed_instr;
  picorv32_axi.picorv32_core.is_lui_auipc_jal <= ff_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal;
  picorv32_axi.picorv32_core.is_lb_lh_lw_lbu_lhu <= ff_buf__picorv32_axi__picorv32_core__is_lb_lh_lw_lbu_lhu;
  picorv32_axi.picorv32_core.is_slli_srli_srai <= ff_buf__picorv32_axi__picorv32_core__is_slli_srli_srai;
  picorv32_axi.picorv32_core.is_jalr_addi_slti_sltiu_xori_ori_andi <= ff_buf__picorv32_axi__picorv32_core__is_jalr_addi_slti_sltiu_xori_ori_andi;
  picorv32_axi.picorv32_core.is_sb_sh_sw <= ff_buf__picorv32_axi__picorv32_core__is_sb_sh_sw;
  picorv32_axi.picorv32_core.is_sll_srl_sra <= ff_buf__picorv32_axi__picorv32_core__is_sll_srl_sra;
  picorv32_axi.picorv32_core.is_lui_auipc_jal_jalr_addi_add_sub <= ff_buf__picorv32_axi__picorv32_core__is_lui_auipc_jal_jalr_addi_add_sub;
  picorv32_axi.picorv32_core.is_slti_blt_slt <= ff_buf__picorv32_axi__picorv32_core__is_slti_blt_slt;
  picorv32_axi.picorv32_core.is_sltiu_bltu_sltu <= ff_buf__picorv32_axi__picorv32_core__is_sltiu_bltu_sltu;
  picorv32_axi.picorv32_core.is_beq_bne_blt_bge_bltu_bgeu <= ff_buf__picorv32_axi__picorv32_core__is_beq_bne_blt_bge_bltu_bgeu;
  picorv32_axi.picorv32_core.is_lbu_lhu_lw <= ff_buf__picorv32_axi__picorv32_core__is_lbu_lhu_lw;
  picorv32_axi.picorv32_core.is_alu_reg_imm <= ff_buf__picorv32_axi__picorv32_core__is_alu_reg_imm;
  picorv32_axi.picorv32_core.is_alu_reg_reg <= ff_buf__picorv32_axi__picorv32_core__is_alu_reg_reg;
  picorv32_axi.picorv32_core.is_compare <= ff_buf__picorv32_axi__picorv32_core__is_compare;
  picorv32_axi.picorv32_core.dbg_rs1val <= ff_buf__picorv32_axi__picorv32_core__dbg_rs1val;
  picorv32_axi.picorv32_core.dbg_rs2val <= ff_buf__picorv32_axi__picorv32_core__dbg_rs2val;
  picorv32_axi.picorv32_core.dbg_rs1val_valid <= ff_buf__picorv32_axi__picorv32_core__dbg_rs1val_valid;
  picorv32_axi.picorv32_core.dbg_rs2val_valid <= ff_buf__picorv32_axi__picorv32_core__dbg_rs2val_valid;
  picorv32_axi.picorv32_core.q_ascii_instr <= ff_buf__picorv32_axi__picorv32_core__q_ascii_instr;
  picorv32_axi.picorv32_core.q_insn_imm <= ff_buf__picorv32_axi__picorv32_core__q_insn_imm;
  picorv32_axi.picorv32_core.q_insn_opcode <= ff_buf__picorv32_axi__picorv32_core__q_insn_opcode;
  picorv32_axi.picorv32_core.q_insn_rs1 <= ff_buf__picorv32_axi__picorv32_core__q_insn_rs1;
  picorv32_axi.picorv32_core.q_insn_rs2 <= ff_buf__picorv32_axi__picorv32_core__q_insn_rs2;
  picorv32_axi.picorv32_core.q_insn_rd <= ff_buf__picorv32_axi__picorv32_core__q_insn_rd;
  picorv32_axi.picorv32_core.dbg_next <= ff_buf__picorv32_axi__picorv32_core__dbg_next;
  picorv32_axi.picorv32_core.dbg_valid_insn <= ff_buf__picorv32_axi__picorv32_core__dbg_valid_insn;
  picorv32_axi.picorv32_core.cached_ascii_instr <= ff_buf__picorv32_axi__picorv32_core__cached_ascii_instr;
  picorv32_axi.picorv32_core.cached_insn_imm <= ff_buf__picorv32_axi__picorv32_core__cached_insn_imm;
  picorv32_axi.picorv32_core.cached_insn_opcode <= ff_buf__picorv32_axi__picorv32_core__cached_insn_opcode;
  picorv32_axi.picorv32_core.cached_insn_rs1 <= ff_buf__picorv32_axi__picorv32_core__cached_insn_rs1;
  picorv32_axi.picorv32_core.cached_insn_rs2 <= ff_buf__picorv32_axi__picorv32_core__cached_insn_rs2;
  picorv32_axi.picorv32_core.cached_insn_rd <= ff_buf__picorv32_axi__picorv32_core__cached_insn_rd;
  picorv32_axi.picorv32_core.cpu_state <= ff_buf__picorv32_axi__picorv32_core__cpu_state;
  picorv32_axi.picorv32_core.irq_state <= ff_buf__picorv32_axi__picorv32_core__irq_state;
  picorv32_axi.picorv32_core.latched_store <= ff_buf__picorv32_axi__picorv32_core__latched_store;
  picorv32_axi.picorv32_core.latched_stalu <= ff_buf__picorv32_axi__picorv32_core__latched_stalu;
  picorv32_axi.picorv32_core.latched_branch <= ff_buf__picorv32_axi__picorv32_core__latched_branch;
  picorv32_axi.picorv32_core.latched_compr <= ff_buf__picorv32_axi__picorv32_core__latched_compr;
  picorv32_axi.picorv32_core.latched_trace <= ff_buf__picorv32_axi__picorv32_core__latched_trace;
  picorv32_axi.picorv32_core.latched_is_lu <= ff_buf__picorv32_axi__picorv32_core__latched_is_lu;
  picorv32_axi.picorv32_core.latched_is_lh <= ff_buf__picorv32_axi__picorv32_core__latched_is_lh;
  picorv32_axi.picorv32_core.latched_is_lb <= ff_buf__picorv32_axi__picorv32_core__latched_is_lb;
  picorv32_axi.picorv32_core.latched_rd <= ff_buf__picorv32_axi__picorv32_core__latched_rd;
  picorv32_axi.picorv32_core.pcpi_timeout_counter <= ff_buf__picorv32_axi__picorv32_core__pcpi_timeout_counter;
  picorv32_axi.picorv32_core.pcpi_timeout <= ff_buf__picorv32_axi__picorv32_core__pcpi_timeout;
  picorv32_axi.picorv32_core.do_waitirq <= ff_buf__picorv32_axi__picorv32_core__do_waitirq;
  picorv32_axi.picorv32_core.alu_out_q <= ff_buf__picorv32_axi__picorv32_core__alu_out_q;
  picorv32_axi.picorv32_core.alu_out_0_q <= ff_buf__picorv32_axi__picorv32_core__alu_out_0_q;
  picorv32_axi.picorv32_core.alu_wait <= ff_buf__picorv32_axi__picorv32_core__alu_wait;
  picorv32_axi.picorv32_core.alu_wait_2 <= ff_buf__picorv32_axi__picorv32_core__alu_wait_2;
  picorv32_axi.picorv32_core.clear_prefetched_high_word_q <= ff_buf__picorv32_axi__picorv32_core__clear_prefetched_high_word_q;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.shift_out <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__shift_out;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.active <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__active;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1 <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2 <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1_q <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs1_q;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2_q <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rs2_q;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd_q <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__rd_q;
  picorv32_axi.picorv32_core.genblk1.pcpi_mul.pcpi_insn_valid_q <= ff_buf__picorv32_axi__picorv32_core__genblk1__pcpi_mul__pcpi_insn_valid_q;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wr_reg <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wr_reg;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_rd_reg <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_rd_reg;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_reg <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_reg;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_ready_reg <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_ready_reg;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_div <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_div;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_divu <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_divu;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_rem <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_rem;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_remu <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__instr_remu;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_q <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__pcpi_wait_q;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.dividend <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__dividend;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.divisor <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__divisor;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient_msk <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__quotient_msk;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.running <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__running;
  picorv32_axi.picorv32_core.genblk2.pcpi_div.outsign <= ff_buf__picorv32_axi__picorv32_core__genblk2__pcpi_div__outsign;
end
// fault injection
always@(posedge inj_flag)begin
  case(inj_id)
    'd0: picorv32_axi.axi_adapter.ack_awvalid <= picorv32_axi.axi_adapter.ack_awvalid^mask[0:0];
    'd1: picorv32_axi.axi_adapter.ack_arvalid <= picorv32_axi.axi_adapter.ack_arvalid^mask[0:0];
    'd2: picorv32_axi.axi_adapter.ack_wvalid <= picorv32_axi.axi_adapter.ack_wvalid^mask[0:0];
    'd3: picorv32_axi.axi_adapter.xfer_done <= picorv32_axi.axi_adapter.xfer_done^mask[0:0];
    'd4: picorv32_axi.picorv32_core.trap_reg <= picorv32_axi.picorv32_core.trap_reg^mask[0:0];
    'd5: picorv32_axi.picorv32_core.mem_valid_reg <= picorv32_axi.picorv32_core.mem_valid_reg^mask[0:0];
    'd6: picorv32_axi.picorv32_core.mem_instr_reg <= picorv32_axi.picorv32_core.mem_instr_reg^mask[0:0];
    'd7: picorv32_axi.picorv32_core.mem_addr_reg <= picorv32_axi.picorv32_core.mem_addr_reg^mask[31:0];
    'd8: picorv32_axi.picorv32_core.mem_wdata_reg <= picorv32_axi.picorv32_core.mem_wdata_reg^mask[31:0];
    'd9: picorv32_axi.picorv32_core.mem_wstrb_reg <= picorv32_axi.picorv32_core.mem_wstrb_reg^mask[3:0];
    'd10: picorv32_axi.picorv32_core.pcpi_valid_reg <= picorv32_axi.picorv32_core.pcpi_valid_reg^mask[0:0];
    'd11: picorv32_axi.picorv32_core.pcpi_insn_reg <= picorv32_axi.picorv32_core.pcpi_insn_reg^mask[31:0];
    'd12: picorv32_axi.picorv32_core.eoi_reg <= picorv32_axi.picorv32_core.eoi_reg^mask[31:0];
    'd13: picorv32_axi.picorv32_core.trace_valid_reg <= picorv32_axi.picorv32_core.trace_valid_reg^mask[0:0];
    'd14: picorv32_axi.picorv32_core.trace_data_reg <= picorv32_axi.picorv32_core.trace_data_reg^mask[35:0];
    'd15: picorv32_axi.picorv32_core.count_cycle <= picorv32_axi.picorv32_core.count_cycle^mask[63:0];
    'd16: picorv32_axi.picorv32_core.count_instr <= picorv32_axi.picorv32_core.count_instr^mask[63:0];
    'd17: picorv32_axi.picorv32_core.reg_pc <= picorv32_axi.picorv32_core.reg_pc^mask[31:0];
    'd18: picorv32_axi.picorv32_core.reg_next_pc <= picorv32_axi.picorv32_core.reg_next_pc^mask[31:0];
    'd19: picorv32_axi.picorv32_core.reg_op1 <= picorv32_axi.picorv32_core.reg_op1^mask[31:0];
    'd20: picorv32_axi.picorv32_core.reg_op2 <= picorv32_axi.picorv32_core.reg_op2^mask[31:0];
    'd21: picorv32_axi.picorv32_core.reg_out <= picorv32_axi.picorv32_core.reg_out^mask[31:0];
    'd22: picorv32_axi.picorv32_core.reg_sh <= picorv32_axi.picorv32_core.reg_sh^mask[4:0];
    'd23: picorv32_axi.picorv32_core.next_insn_opcode <= picorv32_axi.picorv32_core.next_insn_opcode^mask[31:0];
    'd24: picorv32_axi.picorv32_core.dbg_insn_addr <= picorv32_axi.picorv32_core.dbg_insn_addr^mask[31:0];
    'd25: picorv32_axi.picorv32_core.irq_delay <= picorv32_axi.picorv32_core.irq_delay^mask[0:0];
    'd26: picorv32_axi.picorv32_core.irq_active <= picorv32_axi.picorv32_core.irq_active^mask[0:0];
    'd27: picorv32_axi.picorv32_core.irq_mask <= picorv32_axi.picorv32_core.irq_mask^mask[31:0];
    'd28: picorv32_axi.picorv32_core.irq_pending <= picorv32_axi.picorv32_core.irq_pending^mask[31:0];
    'd29: picorv32_axi.picorv32_core.timer <= picorv32_axi.picorv32_core.timer^mask[31:0];
    'd30: picorv32_axi.picorv32_core.cpuregs[0] <= picorv32_axi.picorv32_core.cpuregs[0]^mask[31:0];
    'd31: picorv32_axi.picorv32_core.cpuregs[1] <= picorv32_axi.picorv32_core.cpuregs[1]^mask[31:0];
    'd32: picorv32_axi.picorv32_core.cpuregs[2] <= picorv32_axi.picorv32_core.cpuregs[2]^mask[31:0];
    'd33: picorv32_axi.picorv32_core.cpuregs[3] <= picorv32_axi.picorv32_core.cpuregs[3]^mask[31:0];
    'd34: picorv32_axi.picorv32_core.cpuregs[4] <= picorv32_axi.picorv32_core.cpuregs[4]^mask[31:0];
    'd35: picorv32_axi.picorv32_core.cpuregs[5] <= picorv32_axi.picorv32_core.cpuregs[5]^mask[31:0];
    'd36: picorv32_axi.picorv32_core.cpuregs[6] <= picorv32_axi.picorv32_core.cpuregs[6]^mask[31:0];
    'd37: picorv32_axi.picorv32_core.cpuregs[7] <= picorv32_axi.picorv32_core.cpuregs[7]^mask[31:0];
    'd38: picorv32_axi.picorv32_core.cpuregs[8] <= picorv32_axi.picorv32_core.cpuregs[8]^mask[31:0];
    'd39: picorv32_axi.picorv32_core.cpuregs[9] <= picorv32_axi.picorv32_core.cpuregs[9]^mask[31:0];
    'd40: picorv32_axi.picorv32_core.cpuregs[10] <= picorv32_axi.picorv32_core.cpuregs[10]^mask[31:0];
    'd41: picorv32_axi.picorv32_core.cpuregs[11] <= picorv32_axi.picorv32_core.cpuregs[11]^mask[31:0];
    'd42: picorv32_axi.picorv32_core.cpuregs[12] <= picorv32_axi.picorv32_core.cpuregs[12]^mask[31:0];
    'd43: picorv32_axi.picorv32_core.cpuregs[13] <= picorv32_axi.picorv32_core.cpuregs[13]^mask[31:0];
    'd44: picorv32_axi.picorv32_core.cpuregs[14] <= picorv32_axi.picorv32_core.cpuregs[14]^mask[31:0];
    'd45: picorv32_axi.picorv32_core.cpuregs[15] <= picorv32_axi.picorv32_core.cpuregs[15]^mask[31:0];
    'd46: picorv32_axi.picorv32_core.cpuregs[16] <= picorv32_axi.picorv32_core.cpuregs[16]^mask[31:0];
    'd47: picorv32_axi.picorv32_core.cpuregs[17] <= picorv32_axi.picorv32_core.cpuregs[17]^mask[31:0];
    'd48: picorv32_axi.picorv32_core.cpuregs[18] <= picorv32_axi.picorv32_core.cpuregs[18]^mask[31:0];
    'd49: picorv32_axi.picorv32_core.cpuregs[19] <= picorv32_axi.picorv32_core.cpuregs[19]^mask[31:0];
    'd50: picorv32_axi.picorv32_core.cpuregs[20] <= picorv32_axi.picorv32_core.cpuregs[20]^mask[31:0];
    'd51: picorv32_axi.picorv32_core.cpuregs[21] <= picorv32_axi.picorv32_core.cpuregs[21]^mask[31:0];
    'd52: picorv32_axi.picorv32_core.cpuregs[22] <= picorv32_axi.picorv32_core.cpuregs[22]^mask[31:0];
    'd53: picorv32_axi.picorv32_core.cpuregs[23] <= picorv32_axi.picorv32_core.cpuregs[23]^mask[31:0];
    'd54: picorv32_axi.picorv32_core.cpuregs[24] <= picorv32_axi.picorv32_core.cpuregs[24]^mask[31:0];
    'd55: picorv32_axi.picorv32_core.cpuregs[25] <= picorv32_axi.picorv32_core.cpuregs[25]^mask[31:0];
    'd56: picorv32_axi.picorv32_core.cpuregs[26] <= picorv32_axi.picorv32_core.cpuregs[26]^mask[31:0];
    'd57: picorv32_axi.picorv32_core.cpuregs[27] <= picorv32_axi.picorv32_core.cpuregs[27]^mask[31:0];
    'd58: picorv32_axi.picorv32_core.cpuregs[28] <= picorv32_axi.picorv32_core.cpuregs[28]^mask[31:0];
    'd59: picorv32_axi.picorv32_core.cpuregs[29] <= picorv32_axi.picorv32_core.cpuregs[29]^mask[31:0];
    'd60: picorv32_axi.picorv32_core.cpuregs[30] <= picorv32_axi.picorv32_core.cpuregs[30]^mask[31:0];
    'd61: picorv32_axi.picorv32_core.cpuregs[31] <= picorv32_axi.picorv32_core.cpuregs[31]^mask[31:0];
    'd62: picorv32_axi.picorv32_core.cpuregs[32] <= picorv32_axi.picorv32_core.cpuregs[32]^mask[31:0];
    'd63: picorv32_axi.picorv32_core.cpuregs[33] <= picorv32_axi.picorv32_core.cpuregs[33]^mask[31:0];
    'd64: picorv32_axi.picorv32_core.cpuregs[34] <= picorv32_axi.picorv32_core.cpuregs[34]^mask[31:0];
    'd65: picorv32_axi.picorv32_core.cpuregs[35] <= picorv32_axi.picorv32_core.cpuregs[35]^mask[31:0];
    'd66: picorv32_axi.picorv32_core.mem_state <= picorv32_axi.picorv32_core.mem_state^mask[1:0];
    'd67: picorv32_axi.picorv32_core.mem_wordsize <= picorv32_axi.picorv32_core.mem_wordsize^mask[1:0];
    'd68: picorv32_axi.picorv32_core.mem_rdata_q <= picorv32_axi.picorv32_core.mem_rdata_q^mask[31:0];
    'd69: picorv32_axi.picorv32_core.mem_do_prefetch <= picorv32_axi.picorv32_core.mem_do_prefetch^mask[0:0];
    'd70: picorv32_axi.picorv32_core.mem_do_rinst <= picorv32_axi.picorv32_core.mem_do_rinst^mask[0:0];
    'd71: picorv32_axi.picorv32_core.mem_do_rdata <= picorv32_axi.picorv32_core.mem_do_rdata^mask[0:0];
    'd72: picorv32_axi.picorv32_core.mem_do_wdata <= picorv32_axi.picorv32_core.mem_do_wdata^mask[0:0];
    'd73: picorv32_axi.picorv32_core.mem_la_secondword <= picorv32_axi.picorv32_core.mem_la_secondword^mask[0:0];
    'd74: picorv32_axi.picorv32_core.mem_la_firstword_reg <= picorv32_axi.picorv32_core.mem_la_firstword_reg^mask[0:0];
    'd75: picorv32_axi.picorv32_core.last_mem_valid <= picorv32_axi.picorv32_core.last_mem_valid^mask[0:0];
    'd76: picorv32_axi.picorv32_core.prefetched_high_word <= picorv32_axi.picorv32_core.prefetched_high_word^mask[0:0];
    'd77: picorv32_axi.picorv32_core.mem_16bit_buffer <= picorv32_axi.picorv32_core.mem_16bit_buffer^mask[15:0];
    'd78: picorv32_axi.picorv32_core.instr_lui <= picorv32_axi.picorv32_core.instr_lui^mask[0:0];
    'd79: picorv32_axi.picorv32_core.instr_auipc <= picorv32_axi.picorv32_core.instr_auipc^mask[0:0];
    'd80: picorv32_axi.picorv32_core.instr_jal <= picorv32_axi.picorv32_core.instr_jal^mask[0:0];
    'd81: picorv32_axi.picorv32_core.instr_jalr <= picorv32_axi.picorv32_core.instr_jalr^mask[0:0];
    'd82: picorv32_axi.picorv32_core.instr_beq <= picorv32_axi.picorv32_core.instr_beq^mask[0:0];
    'd83: picorv32_axi.picorv32_core.instr_bne <= picorv32_axi.picorv32_core.instr_bne^mask[0:0];
    'd84: picorv32_axi.picorv32_core.instr_blt <= picorv32_axi.picorv32_core.instr_blt^mask[0:0];
    'd85: picorv32_axi.picorv32_core.instr_bge <= picorv32_axi.picorv32_core.instr_bge^mask[0:0];
    'd86: picorv32_axi.picorv32_core.instr_bltu <= picorv32_axi.picorv32_core.instr_bltu^mask[0:0];
    'd87: picorv32_axi.picorv32_core.instr_bgeu <= picorv32_axi.picorv32_core.instr_bgeu^mask[0:0];
    'd88: picorv32_axi.picorv32_core.instr_lb <= picorv32_axi.picorv32_core.instr_lb^mask[0:0];
    'd89: picorv32_axi.picorv32_core.instr_lh <= picorv32_axi.picorv32_core.instr_lh^mask[0:0];
    'd90: picorv32_axi.picorv32_core.instr_lw <= picorv32_axi.picorv32_core.instr_lw^mask[0:0];
    'd91: picorv32_axi.picorv32_core.instr_lbu <= picorv32_axi.picorv32_core.instr_lbu^mask[0:0];
    'd92: picorv32_axi.picorv32_core.instr_lhu <= picorv32_axi.picorv32_core.instr_lhu^mask[0:0];
    'd93: picorv32_axi.picorv32_core.instr_sb <= picorv32_axi.picorv32_core.instr_sb^mask[0:0];
    'd94: picorv32_axi.picorv32_core.instr_sh <= picorv32_axi.picorv32_core.instr_sh^mask[0:0];
    'd95: picorv32_axi.picorv32_core.instr_sw <= picorv32_axi.picorv32_core.instr_sw^mask[0:0];
    'd96: picorv32_axi.picorv32_core.instr_addi <= picorv32_axi.picorv32_core.instr_addi^mask[0:0];
    'd97: picorv32_axi.picorv32_core.instr_slti <= picorv32_axi.picorv32_core.instr_slti^mask[0:0];
    'd98: picorv32_axi.picorv32_core.instr_sltiu <= picorv32_axi.picorv32_core.instr_sltiu^mask[0:0];
    'd99: picorv32_axi.picorv32_core.instr_xori <= picorv32_axi.picorv32_core.instr_xori^mask[0:0];
    'd100: picorv32_axi.picorv32_core.instr_ori <= picorv32_axi.picorv32_core.instr_ori^mask[0:0];
    'd101: picorv32_axi.picorv32_core.instr_andi <= picorv32_axi.picorv32_core.instr_andi^mask[0:0];
    'd102: picorv32_axi.picorv32_core.instr_slli <= picorv32_axi.picorv32_core.instr_slli^mask[0:0];
    'd103: picorv32_axi.picorv32_core.instr_srli <= picorv32_axi.picorv32_core.instr_srli^mask[0:0];
    'd104: picorv32_axi.picorv32_core.instr_srai <= picorv32_axi.picorv32_core.instr_srai^mask[0:0];
    'd105: picorv32_axi.picorv32_core.instr_add <= picorv32_axi.picorv32_core.instr_add^mask[0:0];
    'd106: picorv32_axi.picorv32_core.instr_sub <= picorv32_axi.picorv32_core.instr_sub^mask[0:0];
    'd107: picorv32_axi.picorv32_core.instr_sll <= picorv32_axi.picorv32_core.instr_sll^mask[0:0];
    'd108: picorv32_axi.picorv32_core.instr_slt <= picorv32_axi.picorv32_core.instr_slt^mask[0:0];
    'd109: picorv32_axi.picorv32_core.instr_sltu <= picorv32_axi.picorv32_core.instr_sltu^mask[0:0];
    'd110: picorv32_axi.picorv32_core.instr_xor <= picorv32_axi.picorv32_core.instr_xor^mask[0:0];
    'd111: picorv32_axi.picorv32_core.instr_srl <= picorv32_axi.picorv32_core.instr_srl^mask[0:0];
    'd112: picorv32_axi.picorv32_core.instr_sra <= picorv32_axi.picorv32_core.instr_sra^mask[0:0];
    'd113: picorv32_axi.picorv32_core.instr_or <= picorv32_axi.picorv32_core.instr_or^mask[0:0];
    'd114: picorv32_axi.picorv32_core.instr_and <= picorv32_axi.picorv32_core.instr_and^mask[0:0];
    'd115: picorv32_axi.picorv32_core.instr_rdcycle <= picorv32_axi.picorv32_core.instr_rdcycle^mask[0:0];
    'd116: picorv32_axi.picorv32_core.instr_rdcycleh <= picorv32_axi.picorv32_core.instr_rdcycleh^mask[0:0];
    'd117: picorv32_axi.picorv32_core.instr_rdinstr <= picorv32_axi.picorv32_core.instr_rdinstr^mask[0:0];
    'd118: picorv32_axi.picorv32_core.instr_rdinstrh <= picorv32_axi.picorv32_core.instr_rdinstrh^mask[0:0];
    'd119: picorv32_axi.picorv32_core.instr_ecall_ebreak <= picorv32_axi.picorv32_core.instr_ecall_ebreak^mask[0:0];
    'd120: picorv32_axi.picorv32_core.instr_fence <= picorv32_axi.picorv32_core.instr_fence^mask[0:0];
    'd121: picorv32_axi.picorv32_core.instr_getq <= picorv32_axi.picorv32_core.instr_getq^mask[0:0];
    'd122: picorv32_axi.picorv32_core.instr_setq <= picorv32_axi.picorv32_core.instr_setq^mask[0:0];
    'd123: picorv32_axi.picorv32_core.instr_retirq <= picorv32_axi.picorv32_core.instr_retirq^mask[0:0];
    'd124: picorv32_axi.picorv32_core.instr_maskirq <= picorv32_axi.picorv32_core.instr_maskirq^mask[0:0];
    'd125: picorv32_axi.picorv32_core.instr_waitirq <= picorv32_axi.picorv32_core.instr_waitirq^mask[0:0];
    'd126: picorv32_axi.picorv32_core.instr_timer <= picorv32_axi.picorv32_core.instr_timer^mask[0:0];
    'd127: picorv32_axi.picorv32_core.decoded_rd <= picorv32_axi.picorv32_core.decoded_rd^mask[5:0];
    'd128: picorv32_axi.picorv32_core.decoded_rs1 <= picorv32_axi.picorv32_core.decoded_rs1^mask[5:0];
    'd129: picorv32_axi.picorv32_core.decoded_rs2 <= picorv32_axi.picorv32_core.decoded_rs2^mask[4:0];
    'd130: picorv32_axi.picorv32_core.decoded_imm <= picorv32_axi.picorv32_core.decoded_imm^mask[31:0];
    'd131: picorv32_axi.picorv32_core.decoded_imm_j <= picorv32_axi.picorv32_core.decoded_imm_j^mask[31:0];
    'd132: picorv32_axi.picorv32_core.decoder_trigger <= picorv32_axi.picorv32_core.decoder_trigger^mask[0:0];
    'd133: picorv32_axi.picorv32_core.decoder_trigger_q <= picorv32_axi.picorv32_core.decoder_trigger_q^mask[0:0];
    'd134: picorv32_axi.picorv32_core.decoder_pseudo_trigger <= picorv32_axi.picorv32_core.decoder_pseudo_trigger^mask[0:0];
    'd135: picorv32_axi.picorv32_core.decoder_pseudo_trigger_q <= picorv32_axi.picorv32_core.decoder_pseudo_trigger_q^mask[0:0];
    'd136: picorv32_axi.picorv32_core.compressed_instr <= picorv32_axi.picorv32_core.compressed_instr^mask[0:0];
    'd137: picorv32_axi.picorv32_core.is_lui_auipc_jal <= picorv32_axi.picorv32_core.is_lui_auipc_jal^mask[0:0];
    'd138: picorv32_axi.picorv32_core.is_lb_lh_lw_lbu_lhu <= picorv32_axi.picorv32_core.is_lb_lh_lw_lbu_lhu^mask[0:0];
    'd139: picorv32_axi.picorv32_core.is_slli_srli_srai <= picorv32_axi.picorv32_core.is_slli_srli_srai^mask[0:0];
    'd140: picorv32_axi.picorv32_core.is_jalr_addi_slti_sltiu_xori_ori_andi <= picorv32_axi.picorv32_core.is_jalr_addi_slti_sltiu_xori_ori_andi^mask[0:0];
    'd141: picorv32_axi.picorv32_core.is_sb_sh_sw <= picorv32_axi.picorv32_core.is_sb_sh_sw^mask[0:0];
    'd142: picorv32_axi.picorv32_core.is_sll_srl_sra <= picorv32_axi.picorv32_core.is_sll_srl_sra^mask[0:0];
    'd143: picorv32_axi.picorv32_core.is_lui_auipc_jal_jalr_addi_add_sub <= picorv32_axi.picorv32_core.is_lui_auipc_jal_jalr_addi_add_sub^mask[0:0];
    'd144: picorv32_axi.picorv32_core.is_slti_blt_slt <= picorv32_axi.picorv32_core.is_slti_blt_slt^mask[0:0];
    'd145: picorv32_axi.picorv32_core.is_sltiu_bltu_sltu <= picorv32_axi.picorv32_core.is_sltiu_bltu_sltu^mask[0:0];
    'd146: picorv32_axi.picorv32_core.is_beq_bne_blt_bge_bltu_bgeu <= picorv32_axi.picorv32_core.is_beq_bne_blt_bge_bltu_bgeu^mask[0:0];
    'd147: picorv32_axi.picorv32_core.is_lbu_lhu_lw <= picorv32_axi.picorv32_core.is_lbu_lhu_lw^mask[0:0];
    'd148: picorv32_axi.picorv32_core.is_alu_reg_imm <= picorv32_axi.picorv32_core.is_alu_reg_imm^mask[0:0];
    'd149: picorv32_axi.picorv32_core.is_alu_reg_reg <= picorv32_axi.picorv32_core.is_alu_reg_reg^mask[0:0];
    'd150: picorv32_axi.picorv32_core.is_compare <= picorv32_axi.picorv32_core.is_compare^mask[0:0];
    'd151: picorv32_axi.picorv32_core.dbg_rs1val <= picorv32_axi.picorv32_core.dbg_rs1val^mask[31:0];
    'd152: picorv32_axi.picorv32_core.dbg_rs2val <= picorv32_axi.picorv32_core.dbg_rs2val^mask[31:0];
    'd153: picorv32_axi.picorv32_core.dbg_rs1val_valid <= picorv32_axi.picorv32_core.dbg_rs1val_valid^mask[0:0];
    'd154: picorv32_axi.picorv32_core.dbg_rs2val_valid <= picorv32_axi.picorv32_core.dbg_rs2val_valid^mask[0:0];
    'd155: picorv32_axi.picorv32_core.q_ascii_instr <= picorv32_axi.picorv32_core.q_ascii_instr^mask[63:0];
    'd156: picorv32_axi.picorv32_core.q_insn_imm <= picorv32_axi.picorv32_core.q_insn_imm^mask[31:0];
    'd157: picorv32_axi.picorv32_core.q_insn_opcode <= picorv32_axi.picorv32_core.q_insn_opcode^mask[31:0];
    'd158: picorv32_axi.picorv32_core.q_insn_rs1 <= picorv32_axi.picorv32_core.q_insn_rs1^mask[4:0];
    'd159: picorv32_axi.picorv32_core.q_insn_rs2 <= picorv32_axi.picorv32_core.q_insn_rs2^mask[4:0];
    'd160: picorv32_axi.picorv32_core.q_insn_rd <= picorv32_axi.picorv32_core.q_insn_rd^mask[4:0];
    'd161: picorv32_axi.picorv32_core.dbg_next <= picorv32_axi.picorv32_core.dbg_next^mask[0:0];
    'd162: picorv32_axi.picorv32_core.dbg_valid_insn <= picorv32_axi.picorv32_core.dbg_valid_insn^mask[0:0];
    'd163: picorv32_axi.picorv32_core.cached_ascii_instr <= picorv32_axi.picorv32_core.cached_ascii_instr^mask[63:0];
    'd164: picorv32_axi.picorv32_core.cached_insn_imm <= picorv32_axi.picorv32_core.cached_insn_imm^mask[31:0];
    'd165: picorv32_axi.picorv32_core.cached_insn_opcode <= picorv32_axi.picorv32_core.cached_insn_opcode^mask[31:0];
    'd166: picorv32_axi.picorv32_core.cached_insn_rs1 <= picorv32_axi.picorv32_core.cached_insn_rs1^mask[4:0];
    'd167: picorv32_axi.picorv32_core.cached_insn_rs2 <= picorv32_axi.picorv32_core.cached_insn_rs2^mask[4:0];
    'd168: picorv32_axi.picorv32_core.cached_insn_rd <= picorv32_axi.picorv32_core.cached_insn_rd^mask[4:0];
    'd169: picorv32_axi.picorv32_core.cpu_state <= picorv32_axi.picorv32_core.cpu_state^mask[7:0];
    'd170: picorv32_axi.picorv32_core.irq_state <= picorv32_axi.picorv32_core.irq_state^mask[1:0];
    'd171: picorv32_axi.picorv32_core.latched_store <= picorv32_axi.picorv32_core.latched_store^mask[0:0];
    'd172: picorv32_axi.picorv32_core.latched_stalu <= picorv32_axi.picorv32_core.latched_stalu^mask[0:0];
    'd173: picorv32_axi.picorv32_core.latched_branch <= picorv32_axi.picorv32_core.latched_branch^mask[0:0];
    'd174: picorv32_axi.picorv32_core.latched_compr <= picorv32_axi.picorv32_core.latched_compr^mask[0:0];
    'd175: picorv32_axi.picorv32_core.latched_trace <= picorv32_axi.picorv32_core.latched_trace^mask[0:0];
    'd176: picorv32_axi.picorv32_core.latched_is_lu <= picorv32_axi.picorv32_core.latched_is_lu^mask[0:0];
    'd177: picorv32_axi.picorv32_core.latched_is_lh <= picorv32_axi.picorv32_core.latched_is_lh^mask[0:0];
    'd178: picorv32_axi.picorv32_core.latched_is_lb <= picorv32_axi.picorv32_core.latched_is_lb^mask[0:0];
    'd179: picorv32_axi.picorv32_core.latched_rd <= picorv32_axi.picorv32_core.latched_rd^mask[5:0];
    'd180: picorv32_axi.picorv32_core.pcpi_timeout_counter <= picorv32_axi.picorv32_core.pcpi_timeout_counter^mask[3:0];
    'd181: picorv32_axi.picorv32_core.pcpi_timeout <= picorv32_axi.picorv32_core.pcpi_timeout^mask[0:0];
    'd182: picorv32_axi.picorv32_core.do_waitirq <= picorv32_axi.picorv32_core.do_waitirq^mask[0:0];
    'd183: picorv32_axi.picorv32_core.alu_out_q <= picorv32_axi.picorv32_core.alu_out_q^mask[31:0];
    'd184: picorv32_axi.picorv32_core.alu_out_0_q <= picorv32_axi.picorv32_core.alu_out_0_q^mask[0:0];
    'd185: picorv32_axi.picorv32_core.alu_wait <= picorv32_axi.picorv32_core.alu_wait^mask[0:0];
    'd186: picorv32_axi.picorv32_core.alu_wait_2 <= picorv32_axi.picorv32_core.alu_wait_2^mask[0:0];
    'd187: picorv32_axi.picorv32_core.clear_prefetched_high_word_q <= picorv32_axi.picorv32_core.clear_prefetched_high_word_q^mask[0:0];
    'd188: picorv32_axi.picorv32_core.genblk1.pcpi_mul.shift_out <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.shift_out^mask[0:0];
    'd189: picorv32_axi.picorv32_core.genblk1.pcpi_mul.active <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.active^mask[3:0];
    'd190: picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1 <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1^mask[32:0];
    'd191: picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2 <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2^mask[32:0];
    'd192: picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1_q <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs1_q^mask[32:0];
    'd193: picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2_q <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.rs2_q^mask[32:0];
    'd194: picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd^mask[63:0];
    'd195: picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd_q <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.rd_q^mask[63:0];
    'd196: picorv32_axi.picorv32_core.genblk1.pcpi_mul.pcpi_insn_valid_q <= picorv32_axi.picorv32_core.genblk1.pcpi_mul.pcpi_insn_valid_q^mask[0:0];
    'd197: picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wr_reg <= picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wr_reg^mask[0:0];
    'd198: picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_rd_reg <= picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_rd_reg^mask[31:0];
    'd199: picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_reg <= picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_reg^mask[0:0];
    'd200: picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_ready_reg <= picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_ready_reg^mask[0:0];
    'd201: picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_div <= picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_div^mask[0:0];
    'd202: picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_divu <= picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_divu^mask[0:0];
    'd203: picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_rem <= picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_rem^mask[0:0];
    'd204: picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_remu <= picorv32_axi.picorv32_core.genblk2.pcpi_div.instr_remu^mask[0:0];
    'd205: picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_q <= picorv32_axi.picorv32_core.genblk2.pcpi_div.pcpi_wait_q^mask[0:0];
    'd206: picorv32_axi.picorv32_core.genblk2.pcpi_div.dividend <= picorv32_axi.picorv32_core.genblk2.pcpi_div.dividend^mask[31:0];
    'd207: picorv32_axi.picorv32_core.genblk2.pcpi_div.divisor <= picorv32_axi.picorv32_core.genblk2.pcpi_div.divisor^mask[62:0];
    'd208: picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient <= picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient^mask[31:0];
    'd209: picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient_msk <= picorv32_axi.picorv32_core.genblk2.pcpi_div.quotient_msk^mask[31:0];
    'd210: picorv32_axi.picorv32_core.genblk2.pcpi_div.running <= picorv32_axi.picorv32_core.genblk2.pcpi_div.running^mask[0:0];
    'd211: picorv32_axi.picorv32_core.genblk2.pcpi_div.outsign <= picorv32_axi.picorv32_core.genblk2.pcpi_div.outsign^mask[0:0];
  endcase
end
// input sequence
always@(posedge tb_clk )begin
  tb_in__resetn <= tb_in2__resetn;
  tb_in__mem_axi_awready <= tb_in2__mem_axi_awready;
  tb_in__mem_axi_wready <= tb_in2__mem_axi_wready;
  tb_in__mem_axi_bvalid <= tb_in2__mem_axi_bvalid;
  tb_in__mem_axi_arready <= tb_in2__mem_axi_arready;
  tb_in__mem_axi_rvalid <= tb_in2__mem_axi_rvalid;
  tb_in__mem_axi_rdata <= tb_in2__mem_axi_rdata;
  tb_in__pcpi_wr <= tb_in2__pcpi_wr;
  tb_in__pcpi_rd <= tb_in2__pcpi_rd;
  tb_in__pcpi_wait <= tb_in2__pcpi_wait;
  tb_in__pcpi_ready <= tb_in2__pcpi_ready;
  tb_in__irq <= tb_in2__irq;
end

endmodule
